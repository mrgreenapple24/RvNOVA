module pc (
    input  wire        clk,
    input  wire        rst,
    input  wire [31:0] pc_next,
    output reg  [31:0] pc
);

    always @(posedge clk or negedge rst) begin
        if (!rst)
            pc <= 32'b0;
        else
            pc <= pc_next;
    end

endmodule
